interface add_if(input logic clk, reset);
    
    logic [7:0] ip1, ip2;
    logic [8:0] out;

endinterface